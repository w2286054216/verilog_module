
/**********************************************************************************************************************************
* File Name:     definition.sv
* Author:          wuqlan
* Email:           
* Date Created:    2022/12/28
* Description:
*
*
* Version:         0.1
*********************************************************************************************************************************/



`ifndef  DEFINITION_SV
`define  DEFINITION_SV

`define  AHB_ADDR_WIDTH    32
`define  AHB_DATA_WIDTH    32

`define  AHB_SLAVE_DEVICES   4

`define  AHB_TRANS_TIMES      40


`endif

