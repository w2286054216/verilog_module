
/**********************************************************************************************************************************
* File Name:     environment.sv
* Author:          wuqlan
* Email:           
* Date Created:    2022/12/28
* Description:      Testbench environment for APB mater interface and APB slave interfaces.
*
*
* Version:         0.1
*********************************************************************************************************************************/


`ifndef  _INCL_ENVIRONMENT
`define  _INCL_ENVIRONMENT

`include "definition.sv"
`include "master_if.sv"
`include "slave_if.sv"
`include "scoreboard.sv"


class Environment;
   
 


endclass


`endif

